library verilog;
use verilog.vl_types.all;
entity cpu_ex is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        iack            : in     vl_logic;
        stall           : in     vl_logic;
        ex_alu_src      : in     vl_logic;
        ex_alu_op       : in     vl_logic_vector(3 downto 0);
        ex_alu_move_cond: in     vl_logic_vector(1 downto 0);
        ex_reg2sn       : in     vl_logic;
        ex_sht          : in     vl_logic;
        ex_shd          : in     vl_logic;
        ex_shp          : in     vl_logic;
        ex_result_sel   : in     vl_logic_vector(1 downto 0);
        ex_reg_dst      : in     vl_logic_vector(1 downto 0);
        ex_memwrite     : in     vl_logic;
        ex_memread      : in     vl_logic;
        ex_store_op     : in     vl_logic_vector(2 downto 0);
        ex_mhi_en       : in     vl_logic;
        ex_mlo_en       : in     vl_logic;
        ex_align_op     : in     vl_logic_vector(2 downto 0);
        ex_mulreg_sel   : in     vl_logic;
        ex_wbdata_sel   : in     vl_logic_vector(1 downto 0);
        ex_regwrite     : in     vl_logic;
        ex_cpwren       : in     vl_logic;
        ex_cprrsel      : in     vl_logic;
        ex_cprrsel      : in     vl_logic;
        ex_w_cp0reg     : in     vl_logic;
        mul_start       : in     vl_logic;
        mul_sign        : in     vl_logic;
        mul_type        : in     vl_logic_vector(1 downto 0);
        wb_regwrite     : in     vl_logic;
        wb_write_num    : in     vl_logic_vector(4 downto 0);
        ex_pca4         : in     vl_logic_vector(31 downto 0);
        ex_ins_rs       : in     vl_logic_vector(4 downto 0);
        ex_ins_rt       : in     vl_logic_vector(4 downto 0);
        ex_ins_rd       : in     vl_logic_vector(4 downto 0);
        ex_ins_sa       : in     vl_logic_vector(4 downto 0);
        ex_a_bus        : in     vl_logic_vector(31 downto 0);
        ex_b_bus        : in     vl_logic_vector(31 downto 0);
        ex_extend_bus   : in     vl_logic_vector(31 downto 0);
        wb_write_bus    : in     vl_logic_vector(31 downto 0);
        mul_a           : in     vl_logic_vector(31 downto 0);
        mul_b           : in     vl_logic_vector(31 downto 0);
        mul_rs          : in     vl_logic_vector(4 downto 0);
        mul_rt          : in     vl_logic_vector(4 downto 0);
        m_memwrite      : out    vl_logic;
        m_memread       : out    vl_logic;
        m_store_op      : out    vl_logic_vector(2 downto 0);
        m_mhi_en        : out    vl_logic;
        m_mlo_en        : out    vl_logic;
        m_align_op      : out    vl_logic_vector(2 downto 0);
        m_mulreg_sel    : out    vl_logic;
        m_wbdata_sel    : out    vl_logic_vector(1 downto 0);
        m_regwrite      : out    vl_logic;
        mul_update_a    : out    vl_logic;
        mul_update_b    : out    vl_logic;
        mul_forward_a   : out    vl_logic_vector(1 downto 0);
        mul_forward_b   : out    vl_logic_vector(1 downto 0);
        mul_stall       : out    vl_logic;
        m_w_cp0reg      : out    vl_logic;
        ex_write_num    : out    vl_logic_vector(4 downto 0);
        m_result_bus    : out    vl_logic_vector(31 downto 0);
        m_b_bus         : out    vl_logic_vector(31 downto 0);
        m_write_num     : out    vl_logic_vector(4 downto 0);
        mul_hi          : out    vl_logic_vector(31 downto 0);
        mul_lo          : out    vl_logic_vector(31 downto 0);
        CPWDBUS         : out    vl_logic_vector(31 downto 0);
        CPWREN          : out    vl_logic;
        CPWRNUM         : out    vl_logic_vector(4 downto 0);
        CPRRNUM         : out    vl_logic_vector(4 downto 0);
        CPRRSEL         : out    vl_logic;
        CPRDBUS         : in     vl_logic_vector(31 downto 0)
    );
end cpu_ex;
