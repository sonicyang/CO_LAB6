library verilog;
use verilog.vl_types.all;
entity fu_shifter_mask is
    port(
        din             : in     vl_logic_vector(4 downto 0);
        dout            : out    vl_logic_vector(31 downto 0)
    );
end fu_shifter_mask;
