library verilog;
use verilog.vl_types.all;
entity forward_unit is
    port(
        ins_rs          : in     vl_logic_vector(4 downto 0);
        ins_rt          : in     vl_logic_vector(4 downto 0);
        m_regwrite      : in     vl_logic;
        m_write_num     : in     vl_logic_vector(4 downto 0);
        wb_regwrite     : in     vl_logic;
        wb_write_num    : in     vl_logic_vector(4 downto 0);
        forward_a       : out    vl_logic_vector(1 downto 0);
        forward_b       : out    vl_logic_vector(1 downto 0)
    );
end forward_unit;
