library verilog;
use verilog.vl_types.all;
entity mul_reg1_ne is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        din             : in     vl_logic;
        wren            : in     vl_logic;
        dout            : out    vl_logic
    );
end mul_reg1_ne;
