library verilog;
use verilog.vl_types.all;
entity mul_fsm is
    generic(
        ST_P1           : integer := 0;
        ST_P2           : integer := 1
    );
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        cs_start        : in     vl_logic;
        phase           : out    vl_logic
    );
end mul_fsm;
