//+FHDR----------------------------------------------------------------
// (C) Copyright CASLab.EE.NCKU
// All Right Reserved
//---------------------------------------------------------------------
// FILE NAME: cpu_decode5to32.v
// AUTHOR: Chen-Chien Wang
// CONTACT INFORMATION: ccwang@casmail.ee.ncku.edu.tw
//---------------------------------------------------------------------
// RELEASE VERSION: V1.0
// VERSION DESCRIPTION: First Edition no errata
//---------------------------------------------------------------------
// RELEASE: 07-27-2004  05:44pm
//---------------------------------------------------------------------
// PURPOSE:
//-FHDR----------------------------------------------------------------

// synopsys translate_off
`include "timescale.v"
// synopsys translate_on

module cpu_decode5to32(din, dout);

        input   [4:0]   din;    // Data input
        output  [31:0]  dout;   // Data Output

        reg     [31:0]  dout;

        always@(din)
        begin

            case(din)
                5'b00000: dout = 32'b00000000000000000000000000000001;
                5'b00001: dout = 32'b00000000000000000000000000000010;
                5'b00010: dout = 32'b00000000000000000000000000000100;
                5'b00011: dout = 32'b00000000000000000000000000001000;
                5'b00100: dout = 32'b00000000000000000000000000010000;
                5'b00101: dout = 32'b00000000000000000000000000100000;
                5'b00110: dout = 32'b00000000000000000000000001000000;
                5'b00111: dout = 32'b00000000000000000000000010000000;
                5'b01000: dout = 32'b00000000000000000000000100000000;
                5'b01001: dout = 32'b00000000000000000000001000000000;
                5'b01010: dout = 32'b00000000000000000000010000000000;
                5'b01011: dout = 32'b00000000000000000000100000000000;
                5'b01100: dout = 32'b00000000000000000001000000000000;
                5'b01101: dout = 32'b00000000000000000010000000000000;
                5'b01110: dout = 32'b00000000000000000100000000000000;
                5'b01111: dout = 32'b00000000000000001000000000000000;
                5'b10000: dout = 32'b00000000000000010000000000000000;
                5'b10001: dout = 32'b00000000000000100000000000000000;
                5'b10010: dout = 32'b00000000000001000000000000000000;
                5'b10011: dout = 32'b00000000000010000000000000000000;
                5'b10100: dout = 32'b00000000000100000000000000000000;
                5'b10101: dout = 32'b00000000001000000000000000000000;
                5'b10110: dout = 32'b00000000010000000000000000000000;
                5'b10111: dout = 32'b00000000100000000000000000000000;
                5'b11000: dout = 32'b00000001000000000000000000000000;
                5'b11001: dout = 32'b00000010000000000000000000000000;
                5'b11010: dout = 32'b00000100000000000000000000000000;
                5'b11011: dout = 32'b00001000000000000000000000000000;
                5'b11100: dout = 32'b00010000000000000000000000000000;
                5'b11101: dout = 32'b00100000000000000000000000000000;
                5'b11110: dout = 32'b01000000000000000000000000000000;
                5'b11111: dout = 32'b10000000000000000000000000000000;

            endcase

        end

endmodule