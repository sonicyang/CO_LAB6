library verilog;
use verilog.vl_types.all;
entity testbench is
    generic(
        CCT             : integer := 10
    );
end testbench;
