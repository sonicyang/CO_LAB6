library verilog;
use verilog.vl_types.all;
entity branch_unit is
    port(
        rs              : in     vl_logic_vector(31 downto 0);
        rt              : in     vl_logic_vector(31 downto 0);
        sel             : in     vl_logic_vector(2 downto 0);
        taken           : out    vl_logic
    );
end branch_unit;
