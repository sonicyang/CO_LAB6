library verilog;
use verilog.vl_types.all;
entity count is
    port(
        go              : in     vl_logic;
        change          : out    vl_logic;
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end count;
